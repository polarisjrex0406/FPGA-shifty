module hex_decoder(input byte x, output byte y);
    // ...
endmodule
