module dec_decoder(input byte x, output byte y);
    assign y = x - 48;
endmodule
